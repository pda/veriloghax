module hello;
  initial
      $display("hello verilog");
endmodule
